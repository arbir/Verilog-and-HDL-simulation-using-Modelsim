module testbench_cmos();
reg t_a,t_b,t_c,t_d,t_e;
wire t_r;
transistor_level innn(t_a,t_b,t_c,t_d,t_e,t_r);
initial begin
	t_a=1'b0;t_b=1'b0;t_c=1'b0;t_d=1'b0;t_e=1'b0;
#1	$display ("The Inputs of Circuit is: a:%d, b:%d, c:%d, d:%d, e:%d ",t_a,t_b,t_c,t_d,t_e );
$display ("The Output of add4 is: %b ",t_r);
#20 t_a=1'b0;t_b=1'b0;t_c=1'b0;t_d=1'b0;t_e=1'b1;
#1	$display ("The Inputs of Circuit is: a:%d, b:%d, c:%d, d:%d, e:%d ",t_a,t_b,t_c,t_d,t_e );
$display ("The Output of add4 is: %b ",t_r);
#20 t_a=1'b0;t_b=1'b0;t_c=1'b0;t_d=1'b1;t_e=1'b0;
#1	$display ("The Inputs of Circuit is: a:%d, b:%d, c:%d, d:%d, e:%d ",t_a,t_b,t_c,t_d,t_e );
$display ("The Output of add4 is: %b ",t_r);
#20 t_a=1'b0;t_b=1'b0;t_c=1'b0;t_d=1'b1;t_e=1'b1;
#1	$display ("The Inputs of Circuit is: a:%d, b:%d, c:%d, d:%d, e:%d ",t_a,t_b,t_c,t_d,t_e );
$display ("The Output of add4 is: %b ",t_r);
#20 t_a=1'b0;t_b=1'b0;t_c=1'b1;t_d=1'b0;t_e=1'b0;
#1	$display ("The Inputs of Circuit is: a:%d, b:%d, c:%d, d:%d, e:%d ",t_a,t_b,t_c,t_d,t_e );
$display ("The Output of add4 is: %b ",t_r);
#20 t_a=1'b0;t_b=1'b0;t_c=1'b1;t_d=1'b0;t_e=1'b1;
#1	$display ("The Inputs of Circuit is: a:%d, b:%d, c:%d, d:%d, e:%d ",t_a,t_b,t_c,t_d,t_e );
$display ("The Output of add4 is: %b ",t_r);
#20 t_a=1'b0;t_b=1'b0;t_c=1'b1;t_d=1'b1;t_e=1'b0;
#1	$display ("The Inputs of Circuit is: a:%d, b:%d, c:%d, d:%d, e:%d ",t_a,t_b,t_c,t_d,t_e );
$display ("The Output of add4 is: %b ",t_r);
#20 t_a=1'b0;t_b=1'b0;t_c=1'b1;t_d=1'b1;t_e=1'b1;
#1	$display ("The Inputs of Circuit is: a:%d, b:%d, c:%d, d:%d, e:%d ",t_a,t_b,t_c,t_d,t_e );
$display ("The Output of add4 is: %b ",t_r);
#20 t_a=1'b0;t_b=1'b1;t_c=1'b0;t_d=1'b0;t_e=1'b0;
#1	$display ("The Inputs of Circuit is: a:%d, b:%d, c:%d, d:%d, e:%d ",t_a,t_b,t_c,t_d,t_e );
$display ("The Output of add4 is: %b ",t_r);
#20 t_a=1'b0;t_b=1'b1;t_c=1'b0;t_d=1'b0;t_e=1'b1;
#1	$display ("The Inputs of Circuit is: a:%d, b:%d, c:%d, d:%d, e:%d ",t_a,t_b,t_c,t_d,t_e );
$display ("The Output of add4 is: %b ",t_r);
#20 t_a=1'b0;t_b=1'b1;t_c=1'b0;t_d=1'b1;t_e=1'b0;
#1	$display ("The Inputs of Circuit is: a:%d, b:%d, c:%d, d:%d, e:%d ",t_a,t_b,t_c,t_d,t_e );
$display ("The Output of add4 is: %b ",t_r);
#20 t_a=1'b0;t_b=1'b1;t_c=1'b0;t_d=1'b1;t_e=1'b1;
#1	$display ("The Inputs of Circuit is: a:%d, b:%d, c:%d, d:%d, e:%d ",t_a,t_b,t_c,t_d,t_e );
$display ("The Output of add4 is: %b ",t_r);
#20 t_a=1'b0;t_b=1'b1;t_c=1'b1;t_d=1'b0;t_e=1'b0;
#1	$display ("The Inputs of Circuit is: a:%d, b:%d, c:%d, d:%d, e:%d ",t_a,t_b,t_c,t_d,t_e );
$display ("The Output of add4 is: %b ",t_r);
#20 t_a=1'b0;t_b=1'b1;t_c=1'b1;t_d=1'b0;t_e=1'b1;
#1	$display ("The Inputs of Circuit is: a:%d, b:%d, c:%d, d:%d, e:%d ",t_a,t_b,t_c,t_d,t_e );
$display ("The Output of add4 is: %b ",t_r);
#20 t_a=1'b0;t_b=1'b1;t_c=1'b1;t_d=1'b1;t_e=1'b0;
#1	$display ("The Inputs of Circuit is: a:%d, b:%d, c:%d, d:%d, e:%d ",t_a,t_b,t_c,t_d,t_e );
$display ("The Output of add4 is: %b ",t_r);
#20 t_a=1'b0;t_b=1'b1;t_c=1'b1;t_d=1'b1;t_e=1'b1;
#1	$display ("The Inputs of Circuit is: a:%d, b:%d, c:%d, d:%d, e:%d ",t_a,t_b,t_c,t_d,t_e );
$display ("The Output of add4 is: %b ",t_r);
#20 t_a=1'b1;t_b=1'b0;t_c=1'b0;t_d=1'b0;t_e=1'b0;
#1	$display ("The Inputs of Circuit is: a:%d, b:%d, c:%d, d:%d, e:%d ",t_a,t_b,t_c,t_d,t_e );
$display ("The Output of add4 is: %b ",t_r);
#20 t_a=1'b1;t_b=1'b0;t_c=1'b0;t_d=1'b0;t_e=1'b1;
#1	$display ("The Inputs of Circuit is: a:%d, b:%d, c:%d, d:%d, e:%d ",t_a,t_b,t_c,t_d,t_e );
$display ("The Output of add4 is: %b ",t_r);
#20 t_a=1'b1;t_b=1'b0;t_c=1'b0;t_d=1'b1;t_e=1'b0;
#1	$display ("The Inputs of Circuit is: a:%d, b:%d, c:%d, d:%d, e:%d ",t_a,t_b,t_c,t_d,t_e );
$display ("The Output of add4 is: %b ",t_r);
#20 t_a=1'b1;t_b=1'b0;t_c=1'b0;t_d=1'b1;t_e=1'b1;
#1	$display ("The Inputs of Circuit is: a:%d, b:%d, c:%d, d:%d, e:%d ",t_a,t_b,t_c,t_d,t_e );
$display ("The Output of add4 is: %b ",t_r);
#20 t_a=1'b1;t_b=1'b0;t_c=1'b1;t_d=1'b0;t_e=1'b0;
#1	$display ("The Inputs of Circuit is: a:%d, b:%d, c:%d, d:%d, e:%d ",t_a,t_b,t_c,t_d,t_e );
$display ("The Output of add4 is: %b ",t_r);
#20 t_a=1'b1;t_b=1'b0;t_c=1'b1;t_d=1'b0;t_e=1'b1;
#1	$display ("The Inputs of Circuit is: a:%d, b:%d, c:%d, d:%d, e:%d ",t_a,t_b,t_c,t_d,t_e );
$display ("The Output of add4 is: %b ",t_r);
#20 t_a=1'b1;t_b=1'b0;t_c=1'b1;t_d=1'b1;t_e=1'b0;
#1	$display ("The Inputs of Circuit is: a:%d, b:%d, c:%d, d:%d, e:%d ",t_a,t_b,t_c,t_d,t_e );
$display ("The Output of add4 is: %b ",t_r);
#20 t_a=1'b1;t_b=1'b0;t_c=1'b1;t_d=1'b1;t_e=1'b1;
#1	$display ("The Inputs of Circuit is: a:%d, b:%d, c:%d, d:%d, e:%d ",t_a,t_b,t_c,t_d,t_e );
$display ("The Output of add4 is: %b ",t_r);
#20 t_a=1'b1;t_b=1'b1;t_c=1'b0;t_d=1'b0;t_e=1'b0;
#1	$display ("The Inputs of Circuit is: a:%d, b:%d, c:%d, d:%d, e:%d ",t_a,t_b,t_c,t_d,t_e );
$display ("The Output of add4 is: %b ",t_r);
#20 t_a=1'b1;t_b=1'b1;t_c=1'b0;t_d=1'b0;t_e=1'b1;
#1	$display ("The Inputs of Circuit is: a:%d, b:%d, c:%d, d:%d, e:%d ",t_a,t_b,t_c,t_d,t_e );
$display ("The Output of add4 is: %b ",t_r);
#20 t_a=1'b1;t_b=1'b1;t_c=1'b0;t_d=1'b1;t_e=1'b0;
#1	$display ("The Inputs of Circuit is: a:%d, b:%d, c:%d, d:%d, e:%d ",t_a,t_b,t_c,t_d,t_e );
$display ("The Output of add4 is: %b ",t_r);
#20 t_a=1'b1;t_b=1'b1;t_c=1'b0;t_d=1'b1;t_e=1'b1;
#1	$display ("The Inputs of Circuit is: a:%d, b:%d, c:%d, d:%d, e:%d ",t_a,t_b,t_c,t_d,t_e );
$display ("The Output of add4 is: %b ",t_r);
#20 t_a=1'b1;t_b=1'b1;t_c=1'b1;t_d=1'b0;t_e=1'b0;
#1	$display ("The Inputs of Circuit is: a:%d, b:%d, c:%d, d:%d, e:%d ",t_a,t_b,t_c,t_d,t_e );
$display ("The Output of add4 is: %b ",t_r);
#20 t_a=1'b1;t_b=1'b1;t_c=1'b1;t_d=1'b0;t_e=1'b1;
#1	$display ("The Inputs of Circuit is: a:%d, b:%d, c:%d, d:%d, e:%d ",t_a,t_b,t_c,t_d,t_e );
$display ("The Output of add4 is: %b ",t_r);
#20 t_a=1'b1;t_b=1'b1;t_c=1'b1;t_d=1'b1;t_e=1'b0;
#1	$display ("The Inputs of Circuit is: a:%d, b:%d, c:%d, d:%d, e:%d ",t_a,t_b,t_c,t_d,t_e );
$display ("The Output of add4 is: %b ",t_r);
#20 t_a=1'b1;t_b=1'b1;t_c=1'b1;t_d=1'b1;t_e=1'b1;
#1	$display ("The Inputs of Circuit is: a:%d, b:%d, c:%d, d:%d, e:%d ",t_a,t_b,t_c,t_d,t_e );
$display ("The Output of add4 is: %b ",t_r);
end
endmodule